netcdf \20120901120000-NCDC-L4_GHRSST-SSTblend-AVHRR_OI-GLOB-v02.0-fv02.0 {
dimensions:
	lat = 720 ;
	lon = 1440 ;
	nv = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float lat(lat) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:axis = "Y" ;
		lat:units = "degrees_north" ;
		lat:valid_min = "-90." ;
		lat:valid_max = "90." ;
		lat:bounds = "lat_bnds" ;
		lat:comment = "uniform grid from -89.875 to 89.875 by 0.25" ;
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:axis = "X" ;
		lon:units = "degrees_east" ;
		lon:valid_min = "-180." ;
		lon:valid_max = "180." ;
		lon:bounds = "lon_bnds" ;
		lon:comment = "uniform grid from -179.875 to 179.875 by 0.25" ;
	int time(time) ;
		time:long_name = "reference time of sst field" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:units = "seconds since 1981-01-01 00:00:00" ;
		time:calendar = "gregorian" ;
		time:comment = "Nominal time because observations are from different sources and are made at different times of the day" ;
	float lat_bnds(lat, nv) ;
		lat_bnds:units = "degress_north" ;
		lat_bnds:comment = "This variable defines the latitude values at the north and south bounds of every 0.25-degree pixel." ;
	float lon_bnds(lon, nv) ;
		lon_bnds:units = "degress_east" ;
		lon_bnds:comment = "This variable defines the longitude values at the west and east bounds of every 0.25-degree pixel." ;
	short analysed_sst(time, lat, lon) ;
		analysed_sst:long_name = "analysed sea surface temperature" ;
		analysed_sst:standard_name = "sea_surface_temperature" ;
		analysed_sst:units = "kelvin" ;
		analysed_sst:_FillValue = -32768s ;
		analysed_sst:add_offset = 273.15f ;
		analysed_sst:scale_factor = 0.01f ;
		analysed_sst:valid_min = -300s ;
		analysed_sst:valid_max = 4500s ;
		analysed_sst:source = "NAVO-L2P-AVHRR19_G, NAVO-L2P-AVHRRMTA_G, NCEP-GTS BUOYS, NCEP-GTS SHIPS, NCEP-ICE50KM" ;
		analysed_sst:comment = "Single-sensor Pathfinder AVHRR SSTs used until 2005; two AVHRRs at a time are used 2006 onward. Sea ice and in situ data used also are ‘near real time’ quality for recent period.  SST (bulk) is at ambiguous depth because multiple types of observations are used." ;
	short analysis_error(time, lat, lon) ;
		analysis_error:long_name = "estimated error standard deviation of analysed_sst" ;
		analysis_error:units = "kelvin" ;
		analysis_error:_FillValue = -32768s ;
		analysis_error:add_offset = 0.f ;
		analysis_error:scale_factor = 0.01f ;
		analysis_error:valid_min = 0s ;
		analysis_error:valid_max = 127s ;
		analysis_error:comment = "Sum of bias, sampling and random errors" ;
	byte mask(time, lat, lon) ;
		mask:long_name = "sea/land field composite mask" ;
		mask:_FillValue = -128b ;
		mask:valid_min = "0b" ;
		mask:valid_max = "1b" ;
		mask:flag_values = "0b,1b" ;
		mask:flag_meanings = "water land" ;
		mask:source = "RWReynolds_landmask_V1.0" ;
		mask:comment = "Binary mask distinguishing water and land only" ;
	byte sea_ice_fraction(time, lat, lon) ;
		sea_ice_fraction:long_name = "sea ice area fraction" ;
		sea_ice_fraction:standard_name = "sea_ice_area_fraction" ;
		sea_ice_fraction:units = "1" ;
		sea_ice_fraction:_FillValue = -128b ;
		sea_ice_fraction:add_offset = 0.f ;
		sea_ice_fraction:scale_factor = 0.01f ;
		sea_ice_fraction:valid_min = 0b ;
		sea_ice_fraction:valid_max = 100b ;
		sea_ice_fraction:source = "NCEP-ICE50KM" ;
		sea_ice_fraction:comment = "7-day median filtered .  Switch from 25 km NASA team ice (http://nsidc.org/data/nsidc-0051.html)  to 50 km NCEP ice (http://polar.ncep.noaa.gov/seaice) after 2004 results in artificial increase in ice coverage." ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:title = "Daily-OI-V2, Final" ;
		:id = "NCDC-L4LRblend-GLOB-AVHRR_OI" ;
		:references = "Reynolds, et al.(2009) What is New in Version 2. Available at http://www.ncdc.noaa.gov/sst/papers/oisst_daily_v02r00_version2-features.pdf;Daily 1/4° Optimum Interpolation Sea Surface Temperature (OISST)- Climate Algorithm Theoretical Theoretical Basis Document, NOAA Climate Data Record Program CDRP-ATBD-0303 Rev. 2 (2013). Available at http://www.ncdc.noaa.gov/cdr/operationalcdrs.html." ;
		:institution = "NOAA/NESDIS/NCDC" ;
		:creator_name = "Viva Banzon" ;
		:creator_email = "viva.banzon@noaa.gov & chunying.liu@noaa.gov" ;
		:creator_url = "http://www.ncdc.noaa.gov/sst/" ;
		:gds_version_id = "v2.0-rev5" ;
		:netcdf_version_id = "4.2.1.1" ;
		:date_created = "2015-07-23" ;
		:product_version = "Version 2.1" ;
		:history = "" ;
		:spatial_resolution = "0.25 degree" ;
		:start_time = "2012-09-01T000000Z" ;
		:stop_time = "2012-09-02T000000Z" ;
		:westernmost_longitude = -179.875f ;
		:easternmost_longitude = 179.875f ;
		:southernmost_latitude = -89.875f ;
		:northernmost_latitude = 89.875f ;
		:file_quality_level = "3" ;
		:source = "NAVO-L2P-AVHRR19_G, NAVO-L2P-AVHRRMTA_G, NCEP-GTS BUOYS, NCEP-GTS SHIPS, NCEP-ICE50KM" ;
		:comment = "WARNING Some applications are unable to properly handle signed byte values. If values are encountered > 127, please subtract 256 from this reported value" ;
		:summary = "NOAA’s ¼-degree Daily Optimum Interpolation Sea Surface temperature (OISST, also known as Reynolds’ SST), currently available as version 2,  is created by interpolating and extrapolating SST observations from different sources, resulting in a smoothed complete field. The sources of data are satellite (AVHRR) and in situ platforms (i.e., ships and buoys), and the specific datasets employed may change over. At the marginal ice zone, sea ice concentrations are used to generate proxy SSTs.  A preliminary version of this file is produced in near-real time (1-day latency), and then replaced with a final version after 2 weeks. Note that this is the AVHRR-ONLY DOISST, available from Oct 1981, but there is a sister DOISST product that includes microwave satellite data, available from June 2002." ;
		:acknowledgement = "This project was supported in part by a grant from the NOAA Climate Data Record (CDR) Program." ;
		:license = "No constraints on data access or use." ;
		:project = "NOAA Optimum Interpolation Sea Surface Temperature (OISST)" ;
		:publisher_name = "OISST Operations Team" ;
		:publisher_email = "oisst_contacts@noaa.gov" ;
		:publisher_url = "http://www.ncdc.noaa.gov/sst" ;
		:naming_authority = "org.ghrsst" ;
		:time_coverage_start = "2012-09-01T000000Z" ;
		:time_coverage_end = "2012-09-02T000000Z" ;
		:platform = "AVHRR-19, MetOpA" ;
		:sensor = "AVHRR_GAC" ;
		:uuid = "46e7d0b7-3bab-4007-9828-c623af70b90f" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "0.25" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "0.25" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:Metadata_Link = "http://doi.org/10.7289/V5SQ8XB5" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory(GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Standard Name Table (v26, 09 November 2012)" ;
		:processing_level = "L4" ;
		:cdm_data_type = "Grid" ;
}
