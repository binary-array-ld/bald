netcdf tmpMwXy8U {
dimensions:
	pdim0 = 11 ;
	pdim1 = 17 ;
variables:
	int parent_variable(pdim0, pdim1) ;
		parent_variable:rdf__type = "bald__Array" ;
		parent_variable:SDN_ParameterDiscoveryCode = "BactTaxaAbundSed" ;
		parent_variable:submursible_name = "Nautilus" ;

	int prefix_list ;
		prefix_list:bald__ = "http://binary-array-ld.net/latest/" ;
		prefix_list:rdf__ = "http://www.w3.org/1999/02/22-rdf-syntax-ns#" ;

	int alias_list ;
		alias_list:SDN_ParameterDiscoveryCode = "http://vocab.nerc.ac.uk/isoCodelists/sdnCodelists/cdicsrCodeList.xml#SDN_ParameterDiscoveryCode" ;
		alias_list:BactTaxaAbundSed = "http://vocab.nerc.ac.uk/collection/P02/current/BAUC/" ;


// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:rdf__type = "bald__Container" ;
		:bald__isPrefixedBy = "prefix_list" ;
		:bald__isAliasedBy = "alias_list" ;

}
