netcdf tmpMwXy8U {
dimensions:
	pdim0 = 11 ;
	pdim1 = 17 ;
variables:
        int prefix_list(pdim0, pdim1) ;
  		prefix_list:bald__ = "http://binary-array-ld.net/latest/" ;
		prefix_list:metce__ = "http://codes.wmo.int/common/observation-type/METCE/2013/" ;
  		prefix_list:rdf__ = "http://www.w3.org/1999/02/22-rdf-syntax-ns#" ;
		
	int data_variable1(pdim0, pdim1) ;
		data_variable1:bald__references = "location_variable" ;
		data_variable1:long_name = "Gerald";
		data_variable1:obtype = "metce__SamplingObservation";

        int data_variable2(pdim0, pdim1) ;
		data_variable2:bald__references = "location_variable" ;
		data_variable2:long_name = "Imelda";
		data_variable2:obtype = "metce__SamplingObservation";

        int pdim0(pdim0) ;

        int pdim1(pdim1) ;

	int location_variable(pdim0, pdim1) ;
	        location_variable:rdf__type = "bald__Reference";
		location_variable:bald__array = "location_variable" ;
		location_variable:bald__references = "location_reference_system" ;

	int location_reference_system;
	        location_variable:rdf__type = "bald__Reference";
	        location_reference_system:bald__array = "location_reference_system";
		location_reference_system:pcode = "4897";

	int set_collection ;
	        set_collection:bald__references = "data_variable1 data_variable2" ;

	int list_collection ;
	        list_collection:bald__references = "data_variable1,data_variable2" ;


// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:bald__isPrefixedBy = "prefix_list" ;

}
