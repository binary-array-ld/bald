netcdf GEMS_CO2_Apr2006 {
dimensions:
	longitude = 360 ;
	latitude = 181 ;
	levelist = 60 ;
	time = 1 ;
variables:
	float longitude(longitude) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	float latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	int levelist(levelist) ;
		levelist:long_name = "model_level_number" ;
	int time(time) ;
		time:units = "hours since 1900-01-01 00:00:0.0" ;
		time:standard_name = "time" ;
	short co2(time, levelist, latitude, longitude) ;
		co2:scale_factor = 0.000981685145029486 ;
		co2:add_offset = 403.192219379918 ;
		co2:_FillValue = -32767s ;
		co2:missing_value = -32767s ;
		co2:units = "kg kg**-1" ;
		co2:long_name = "Carbon Dioxide" ;
		co2:standard_name = "mass_fraction_of_carbon_dioxide_in_air" ;
	short lnsp(time, levelist, latitude, longitude) ;
		lnsp:scale_factor = 1.03952457840347e-05 ;
		lnsp:add_offset = 11.2087164280841 ;
		lnsp:_FillValue = -32767s ;
		lnsp:missing_value = -32767s ;
		lnsp:long_name = "Logarithm of surface pressure" ;

// global attributes:
		:Conventions = "CF-1.0" ;

data:

 longitude = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 
    190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 
    204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 
    218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 
    232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 
    246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 
    260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 
    274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 
    288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 
    302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 
    316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 
    330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 
    344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 
    358, 359 ;

 latitude = 90, 89, 88, 87, 86, 85, 84, 83, 82, 81, 80, 79, 78, 77, 76, 75, 
    74, 73, 72, 71, 70, 69, 68, 67, 66, 65, 64, 63, 62, 61, 60, 59, 58, 57, 
    56, 55, 54, 53, 52, 51, 50, 49, 48, 47, 46, 45, 44, 43, 42, 41, 40, 39, 
    38, 37, 36, 35, 34, 33, 32, 31, 30, 29, 28, 27, 26, 25, 24, 23, 22, 21, 
    20, 19, 18, 17, 16, 15, 14, 13, 12, 11, 10, 9, 8, 7, 6, 5, 4, 3, 2, 1, 0, 
    -1, -2, -3, -4, -5, -6, -7, -8, -9, -10, -11, -12, -13, -14, -15, -16, 
    -17, -18, -19, -20, -21, -22, -23, -24, -25, -26, -27, -28, -29, -30, 
    -31, -32, -33, -34, -35, -36, -37, -38, -39, -40, -41, -42, -43, -44, 
    -45, -46, -47, -48, -49, -50, -51, -52, -53, -54, -55, -56, -57, -58, 
    -59, -60, -61, -62, -63, -64, -65, -66, -67, -68, -69, -70, -71, -72, 
    -73, -74, -75, -76, -77, -78, -79, -80, -81, -82, -83, -84, -85, -86, 
    -87, -88, -89, -90 ;

 levelist = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60 ;

 time = 931344 ;
}
