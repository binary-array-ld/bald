netcdf tmpMwXy8U {
dimensions:
	pdim0 = 11 ;
	pdim1 = 17 ;
variables:
	int parent_variable(pdim0, pdim1) ;
		parent_variable:rdf__type = "bald__Array" ;
		parent_variable:bald__references = "child_variable" ;
	int child_variable(pdim0, pdim1) ;
		child_variable:rdf__type = "bald__Reference" ;
		child_variable:bald__array = "child_variable" ;
	int prefix_list ;
		prefix_list:bald__ = "http://binary-array-ld.net/latest/" ;
		prefix_list:rdf__ = "http://www.w3.org/1999/02/22-rdf-syntax-ns#" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:rdf__type = "bald__Container" ;
		:bald__isPrefixedBy = "prefix_list" ;
}
