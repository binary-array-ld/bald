netcdf tmpMwXy8U {
dimensions:
        x_t = 144 ;
	y_t = 91 ;
        x_q = 144 ;
	y_q = 90 ;
	time = 4 ;
variables:
        float x_t(x_t) ;
	    x_t:cf__standard_name = "longitude" ;
	    x_t:nc__units = "degrees" ;


	float y_t(y_t) ;
	    y_t:cf__standard_name = "latitude" ;
	    y_t:nc__units = "degrees" ;


        float x_q(x_q) ;
	    x_q:cf__standard_name = "longitude" ;
	    x_q:nc__units = "degrees" ;


	float y_q(y_q) ;
	    y_q:cf__standard_name = "latitude" ;
	    y_q:nc__units = "degrees" ;

        int theta_points ;
	    theta_points:georef__wkt_crs = "http://www.epsg-registry.org/export.htm?wkt=urn:ogc:def:crs:EPSG::4326" ;
	    theta_points:georef__coord_tuple = "(y_t x_t)" ;
	    theta_points:rdfs__label = "Theta Points" ;
	    theta_points:dct__description = "Arakawa C Theta points defined with respect to a 2D WGS84 geodetic surface." ;

        int u_points ;
	    u_points:cf__wkt_crs = "http://www.epsg-registry.org/export.htm?wkt=urn:ogc:def:crs:EPSG::4326" ;
	    u_points:georef__coord_tuple = "(y_t x_q)" ;
	    u_points:rdfs__label = "U Points" ;
	    u_points:dct__description = "Arakawa C U points defined with respect to a 2D WGS84 geodetic surface." ;

        int v_points ;
	    v_points:georef__wkt_crs = "http://www.epsg-registry.org/export.htm?wkt=urn:ogc:def:crs:EPSG::4326" ;
	    v_points:georef__coord_tuple = "(y_q x_t)" ;
	    v_points:rdfs__label = "V Points" ;
	    v_points:dct__description = "Arakawa C V points defined with respect to a 2D WGS84 geodetic surface." ;

	string time(time) ;
	    time:rdfs__label = "Time" ;

// global attributes:
		:bald__isPrefixedBy = "prefix_list" ;

data:

y_t = -90, -88, -86, -84, -82, -80, -78, -76, -74, -72, -70, -68, -66, -64, -62, -60, -58, -56, -54, -52, -50, -48, -46, -44, -42, -40, -38, -36, -34, -32, -30, -28, -26, -24, -22, -20, -18, -16, -14, -12, -10, -8, -6, -4, -2, 0, 2, 4, 6, 8, 10, 12, 14, 16, 18, 20, 22, 24, 26, 28, 30, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 62, 64, 66, 68, 70, 72, 74, 76, 78, 80, 82, 84, 86, 88, 90 ;

x_t = 0.0, 2.5, 5.0, 7.5, 10.0, 12.5, 15.0, 17.5, 20.0, 22.5, 25.0, 27.5, 30.0, 32.5, 35.0, 37.5, 40.0, 42.5, 45.0, 47.5, 50.0, 52.5, 55.0, 57.5, 60.0, 62.5, 65.0, 67.5, 70.0, 72.5, 75.0, 77.5, 80.0, 82.5, 85.0, 87.5, 90.0, 92.5, 95.0, 97.5, 100.0, 102.5, 105.0, 107.5, 110.0, 112.5, 115.0, 117.5, 120.0, 122.5, 125.0, 127.5, 130.0, 132.5, 135.0, 137.5, 140.0, 142.5, 145.0, 147.5, 150.0, 152.5, 155.0, 157.5, 160.0, 162.5, 165.0, 167.5, 170.0, 172.5, 175.0, 177.5, 180.0, 182.5, 185.0, 187.5, 190.0, 192.5, 195.0, 197.5, 200.0, 202.5, 205.0, 207.5, 210.0, 212.5, 215.0, 217.5, 220.0, 222.5, 225.0, 227.5, 230.0, 232.5, 235.0, 237.5, 240.0, 242.5, 245.0, 247.5, 250.0, 252.5, 255.0, 257.5, 260.0, 262.5, 265.0, 267.5, 270.0, 272.5, 275.0, 277.5, 280.0, 282.5, 285.0, 287.5, 290.0, 292.5, 295.0, 297.5, 300.0, 302.5, 305.0, 307.5, 310.0, 312.5, 315.0, 317.5, 320.0, 322.5, 325.0, 327.5, 330.0, 332.5, 335.0, 337.5, 340.0, 342.5, 345.0, 347.5, 350.0, 352.5, 355.0, 357.5 ;

y_q = -89, -87, -85, -83, -81, -79, -77, -75, -73, -71, -69, -67, -65, -63, -61, -59, -57, -55, -53, -51, -49, -47, -45, -43, -41, -39, -37, -35, -33, -31, -29, -27, -25, -23, -21, -19, -17, -15, -13, -11, -9, -7, -5, -3, -1, 1, 3, 5, 7, 9, 11, 13, 15, 17, 19, 21, 23, 25, 27, 29, 31, 33, 35, 37, 39, 41, 43, 45, 47, 49, 51, 53, 55, 57, 59, 61, 63, 65, 67, 69, 71, 73, 75, 77, 79, 81, 83, 85, 87, 89 ;

x_q = 1.25, 3.75, 6.25, 8.75, 11.25, 13.75, 16.25, 18.75, 21.25, 23.75, 26.25, 28.75, 31.25, 33.75, 36.25, 38.75, 41.25, 43.75, 46.25, 48.75, 51.25, 53.75, 56.25, 58.75, 61.25, 63.75, 66.25, 68.75, 71.25, 73.75, 76.25, 78.75, 81.25, 83.75, 86.25, 88.75, 91.25, 93.75, 96.25, 98.75, 101.25, 103.75, 106.25, 108.75, 111.25, 113.75, 116.25, 118.75, 121.25, 123.75, 126.25, 128.75, 131.25, 133.75, 136.25, 138.75, 141.25, 143.75, 146.25, 148.75, 151.25, 153.75, 156.25, 158.75, 161.25, 163.75, 166.25, 168.75, 171.25, 173.75, 176.25, 178.75, 181.25, 183.75, 186.25, 188.75, 191.25, 193.75, 196.25, 198.75, 201.25, 203.75, 206.25, 208.75, 211.25, 213.75, 216.25, 218.75, 221.25, 223.75, 226.25, 228.75, 231.25, 233.75, 236.25, 238.75, 241.25, 243.75, 246.25, 248.75, 251.25, 253.75, 256.25, 258.75, 261.25, 263.75, 266.25, 268.75, 271.25, 273.75, 276.25, 278.75, 281.25, 283.75, 286.25, 288.75, 291.25, 293.75, 296.25, 298.75, 301.25, 303.75, 306.25, 308.75, 311.25, 313.75, 316.25, 318.75, 321.25, 323.75, 326.25, 328.75, 331.25, 333.75, 336.25, 338.75, 341.25, 343.75, 346.25, 348.75, 351.25, 353.75, 356.25, 358.75 ;

time = "2020-05-05T00:00Z", "2020-05-05T06:00Z", "2020-05-05T12:00Z", "2020-05-05T18:00Z" ;

// prefix group
group: prefix_list {
    :bald__ = "https://www.opengis.net/def/binary-array-ld/" ;
    :rdf__ = "http://www.w3.org/1999/02/22-rdf-syntax-ns#" ;
    :bald__ = "https://www.opengis.net/def/binary-array-ld/" ;
    :rdf__ = "http://www.w3.org/1999/02/22-rdf-syntax-ns#" ;
    :rdfs__ = "http://www.w3.org/2000/01/rdf-schema#" ;
    :cf__ = "http://def.scitools.org.uk/CFTerms/" ;
    :nc__ = "http://def.scitools.org.uk/NetCDF/" ;
    :geo__ = "http://www.opengis.net/ont/geosparql#" ;
    :nc__ = "http://def.scitools.org.uk/NetCDF/" ;
    :georef__ = "http://def.scitools.org.uk/referencing-by-coordinates/" ;
    :dct__ = "http://purl.org/dc/terms/" ;
}

group: vector_quantities {
    :vq__vector_quantities = "wind" ;


group: wind {
variables:

    float u_wind(time, y_t, x_q) ;
        u_wind:cf__standard_name = "x_wind" ;
	u_wind:nc__units = "m s-1" ;
        u_wind:georef__domain = "u_points" ;

    float v_wind(time, y_q, x_t) ;
        v_wind:cf__standard_name = "y_wind" ;
	v_wind:nc__units = "m s-1" ;
        v_wind:georef__domain = "v_points" ;

    :vq__i_component = "x_wind" ;
    :vq__j_component = "y_wind" ;
    :rdfs__label = "Wind Vector" ;
}

}

group: scalar_quantities {
variables:

    float air_pressure(time, y_t, x_t) ;
        air_pressure:cf__standard_name = "air_pressure" ;
	air_pressure:nc__units = "Pa" ;
	air_pressure:georef__domain = "theta_points" ;

}

}
