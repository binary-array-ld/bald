netcdf tmpcdltest {
variables:
        int gfsmos_process_chain;
        gfsmos_process_chain:OM_Process = "(step1 step2)";

int step1;
        step1:LE_ProcessStep = "NWP__/Models/GFS13" ;
        step1:LE_Source = "DA__/Methods/GDAS13" ;

int step2 ;
        step2:LE_ProcessStep = "StatPP__/Methods/GFSMOS05" ;
        step2:LE_Source = "NWP__/Models/GFS13" ;

//global attribute
        :process_chain = "gfsmos_process_chain";
        :bald__isPrefixedBy = "prefix_list" ;

group: prefix_list {

// group attributes:
        :DA = "https://codes.nws.noaa.gov/DataAssimilation" ;
        :NWP = "https://codes.nws.noaa.gov/NumericalWeatherPrediction" ;
        :StatPP = "https://codes.nws.noaa.gov/StatisticalPostProcessing" ;
        :bald = "http://binary-array-ld.net/latest/" ;
      
  } // group bald__prefix_list
}
