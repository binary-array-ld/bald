netcdf trajectory_AfricanEasterlyWave {
dimensions:
	trajectory = 493 ;
	sample = 10732 ;
variables:
	int count(trajectory) ;
		count:long_name = "number of observations for the easterly wave" ;
		count:sample_dimension = "sample" ;
	int trajectory(trajectory) ;
		trajectory:long_name = "easterly wave trajectory" ;
		trajectory:cf_role = "trajectory_id" ;
	float time(sample) ;
		time:_FillValue = -999.f ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "days since 1900-01-01 00:00:00" ;
		time:calendar = "gregorian" ;
		time:axis = "T" ;
	float lat(sample) ;
		lat:_FillValue = -999.f ;
		lat:long_name = "wave trough centroid latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:cell_methods = "latitude: mean (over the wave trough)" ;
	float lon(sample) ;
		lon:_FillValue = -999.f ;
		lon:long_name = "wave trough centroid longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:cell_methods = "longitude: mean (over the wave trough)" ;
	float maxlat(sample) ;
		maxlat:_FillValue = -999.f ;
		maxlat:long_name = "wave trough maximum latitude" ;
		maxlat:units = "degrees_north" ;
		maxlat:coordinates = "time lat lon" ;
		maxlat:cell_methods = "latitude: maximum (over the wave trough)" ;
	float meanlonatmaxlat(sample) ;
		meanlonatmaxlat:_FillValue = -999.f ;
		meanlonatmaxlat:long_name = "mean longitude of wave trough maximum latitude" ;
		meanlonatmaxlat:units = "degrees_east" ;
		meanlonatmaxlat:coordinates = "time lat lon" ;
		meanlonatmaxlat:cell_methods = "latitude: maximum (over the wave trough) longitude: mean (across the wave trough at maximum latitude)" ;
	float minlat(sample) ;
		minlat:_FillValue = -999.f ;
		minlat:long_name = "wave trough minimum latitude" ;
		minlat:units = "degrees_north" ;
		minlat:coordinates = "time lat lon" ;
		minlat:cell_methods = "latitude: minimum (over the wave trough)" ;
	float meanlonatminlat(sample) ;
		meanlonatminlat:_FillValue = -999.f ;
		meanlonatminlat:long_name = "mean longitude of wave trough minimum latitude" ;
		meanlonatminlat:units = "degrees_east" ;
		meanlonatminlat:coordinates = "time lat lon" ;
		meanlonatminlat:cell_methods = "latitude: minimum (over the wave trough) longitude: mean (across the wave trough at minimum latitude)" ;
	float wavelength(sample) ;
		wavelength:_FillValue = -999.f ;
		wavelength:long_name = "horizontal wavelength" ;
		wavelength:units = "km" ;
		wavelength:coordinates = "time lat lon" ;
		wavelength:comment = "wavelength defined as distance in wave direction where curvature vorticity anomaly for wave trough equals 0 s-1." ;
	float meanrv(sample) ;
		meanrv:_FillValue = -999.f ;
		meanrv:long_name = "wave trough mean relative vorticity" ;
		meanrv:units = "s-1" ;
		meanrv:coordinates = "time lat lon" ;
		meanrv:cell_methods = "area: mean (over the wave trough)" ;
	float maxrv(sample) ;
		maxrv:_FillValue = -999.f ;
		maxrv:long_name = "wave trough maximum relative vorticity" ;
		maxrv:units = "s-1" ;
		maxrv:coordinates = "time lat lon" ;
		maxrv:cell_methods = "area: maximum (over the wave trough)" ;
	float minrv(sample) ;
		minrv:_FillValue = -999.f ;
		minrv:long_name = "wave trough minimum relative vorticity" ;
		minrv:units = "s-1" ;
		minrv:coordinates = "time lat lon" ;
		minrv:cell_methods = "area: minimum (over the wave trough)" ;
	float stdrv(sample) ;
		stdrv:_FillValue = -999.f ;
		stdrv:long_name = "wave trough standard deviation relative vorticity" ;
		stdrv:units = "s-1" ;
		stdrv:coordinates = "time lat lon" ;
		stdrv:cell_methods = "area: standard_deviation (over the wave trough)" ;
	float meancrv(sample) ;
		meancrv:_FillValue = -999.f ;
		meancrv:long_name = "wave trough mean curvature vorticity" ;
		meancrv:units = "s-1" ;
		meancrv:coordinates = "time lat lon" ;
		meancrv:cell_methods = "area: mean (over the wave trough)" ;
	float maxcrv(sample) ;
		maxcrv:_FillValue = -999.f ;
		maxcrv:long_name = "wave trough maximum curvature vorticity" ;
		maxcrv:units = "s-1" ;
		maxcrv:coordinates = "time lat lon" ;
		maxcrv:cell_methods = "area: maximum (over the wave trough)" ;
	float mincrv(sample) ;
		mincrv:_FillValue = -999.f ;
		mincrv:long_name = "wave trough minimum curvature vorticity" ;
		mincrv:units = "s-1" ;
		mincrv:coordinates = "time lat lon" ;
		mincrv:cell_methods = "area: minimum (over the wave trough)" ;
	float stdcrv(sample) ;
		stdcrv:_FillValue = -999.f ;
		stdcrv:long_name = "wave trough standard deviation curvature vorticity" ;
		stdcrv:units = "s-1" ;
		stdcrv:coordinates = "time lat lon" ;
		stdcrv:cell_methods = "area: standard_deviation (over the wave trough)" ;
	float meansrv(sample) ;
		meansrv:_FillValue = -999.f ;
		meansrv:long_name = "wave trough mean shear vorticity" ;
		meansrv:units = "s-1" ;
		meansrv:coordinates = "time lat lon" ;
		meansrv:cell_methods = "area: mean (over the wave trough)" ;
	float maxsrv(sample) ;
		maxsrv:_FillValue = -999.f ;
		maxsrv:long_name = "wave trough maximum shear vorticity" ;
		maxsrv:units = "s-1" ;
		maxsrv:coordinates = "time lat lon" ;
		maxsrv:cell_methods = "area: maximum (over the wave trough)" ;
	float minsrv(sample) ;
		minsrv:_FillValue = -999.f ;
		minsrv:long_name = "wave trough minimum shear vorticity" ;
		minsrv:units = "s-1" ;
		minsrv:coordinates = "time lat lon" ;
		minsrv:cell_methods = "area: minimum (over the wave trough)" ;
	float stdsrv(sample) ;
		stdsrv:_FillValue = -999.f ;
		stdsrv:long_name = "wave trough standard deviation shear vorticity" ;
		stdsrv:units = "s-1" ;
		stdsrv:coordinates = "time lat lon" ;
		stdsrv:cell_methods = "area: standard_deviation (over the wave trough)" ;
	float meanolr(sample) ;
		meanolr:_FillValue = -999.f ;
		meanolr:long_name = "wave trough mean outgoing longwave radiation" ;
		meanolr:units = "W m-2" ;
		meanolr:coordinates = "time lat lon" ;
		meanolr:cell_methods = "area: mean (over the wave trough)" ;
		meanolr:source = "The Outgoing Longwave Radiation - Daily CDR used in this study was acquired from NOAA\'s National Climatic Data Center (http://www.ncdc.noaa.gov).  This CDR was originally developed by Hai-Tien Lee and colleagues for the NOAA\'s CDR Program." ;
		meanolr:references = "Lee,H.-T., C.J. Schreck, K. R. Knapp, 2014: Generation of the Daily OLR Climate Data Record.  2014 EUMETSTAT Meteorological Satellite Conference, 22-26 September 2014, Geneva, Switzerland." ;
	float stdolr(sample) ;
		stdolr:_FillValue = -999.f ;
		stdolr:long_name = "wave trough standard deviation outgoing longwave radiation" ;
		stdolr:units = "W m-2" ;
		stdolr:coordinates = "time lat lon" ;
		stdolr:cell_methods = "area: standard_deviation (over the wave trough)" ;
		stdolr:source = "The Outgoing Longwave Radiation - Daily CDR used in this study was acquired from NOAA\'s National Climatic Data Center (http://www.ncdc.noaa.gov).  This CDR was originally developed by Hai-Tien Lee and colleagues for the NOAA\'s CDR Program." ;
		stdolr:references = "Lee,H.-T., C.J. Schreck, K. R. Knapp, 2014: Generation of the Daily OLR Climate Data Record.  2014 EUMETSTAT Meteorological Satellite Conference, 22-26 September 2014, Geneva, Switzerland." ;
	float olr_area_fraction(sample) ;
		olr_area_fraction:_FillValue = -999.f ;
		olr_area_fraction:long_name = "wave trough outgoing longwave radiation area fraction" ;
		olr_area_fraction:units = "" ;
		olr_area_fraction:coordinates = "time lat lon" ;
		olr_area_fraction:source = "The Outgoing Longwave Radiation - Daily CDR used in this study was acquired from NOAA\'s National Climatic Data Center (http://www.ncdc.noaa.gov).  This CDR was originally developed by Hai-Tien Lee and colleagues for the NOAA\'s CDR Program." ;
		olr_area_fraction:references = "Lee,H.-T., C.J. Schreck, K. R. Knapp, 2014: Generation of the Daily OLR Climate Data Record.  2014 EUMETSTAT Meteorological Satellite Conference, 22-26 September 2014, Geneva, Switzerland." ;
		olr_area_fraction:comment = "Fractional area coverage of available OLR data for the wave trough." ;
	float meanolra(sample) ;
		meanolra:_FillValue = -999.f ;
		meanolra:long_name = "wave trough mean outgoing longwave radiation anomalies" ;
		meanolra:units = "W m-2" ;
		meanolra:coordinates = "time lat lon" ;
		meanolra:cell_methods = "area: mean (over the wave trough)" ;
		meanolra:source = "The Outgoing Longwave Radiation - Daily CDR used in this study was acquired from NOAA\'s National Climatic Data Center (http://www.ncdc.noaa.gov).  This CDR was originally developed by Hai-Tien Lee and colleagues for the NOAA\'s CDR Program." ;
		meanolra:references = "Lee,H.-T., C.J. Schreck, K. R. Knapp, 2014: Generation of the Daily OLR Climate Data Record.  2014 EUMETSTAT Meteorological Satellite Conference, 22-26 September 2014, Geneva, Switzerland." ;
		meanolra:comment = "OLR anomalies calculated by removing daily OLR from the long-term daily mean for 1981-2010." ;
	float stdolra(sample) ;
		stdolra:_FillValue = -999.f ;
		stdolra:long_name = "wave trough standard deviation outgoing longwave radiation anomalies" ;
		stdolra:units = "W m-2" ;
		stdolra:coordinates = "time lat lon" ;
		stdolra:cell_methods = "area: standard_deviation (over the wave trough)" ;
		stdolra:source = "The Outgoing Longwave Radiation - Daily CDR used in this study was acquired from NOAA\'s National Climatic Data Center (http://www.ncdc.noaa.gov).  This CDR was originally developed by Hai-Tien Lee and colleagues for the NOAA\'s CDR Program." ;
		stdolra:references = "Lee,H.-T., C.J. Schreck, K. R. Knapp, 2014: Generation of the Daily OLR Climate Data Record.  2014 EUMETSTAT Meteorological Satellite Conference, 22-26 September 2014, Geneva, Switzerland." ;
		stdolra:comment = "OLR anomalies calculated by removing daily OLR from the long-term daily mean for 1981-2010." ;
	float meanctb(sample) ;
		meanctb:_FillValue = -999.f ;
		meanctb:long_name = "wave trough mean Claus brightness temperature" ;
		meanctb:units = "K" ;
		meanctb:coordinates = "time lat lon" ;
		meanctb:cell_methods = "area: mean (over the wave trough)" ;
		meanctb:references = "Environmental Systems Science Centre (ESSC), [Robinson, G.J.] . Cloud Archive User Service (CLAUS), [Internet]. NCAS British Atmospheric Data Centre, 2002. Available from http://badc.nerc.ac.uk/view/badc.nerc.ac.uk__ATOM__dataent_claus." ;
	float stdctb(sample) ;
		stdctb:_FillValue = -999.f ;
		stdctb:long_name = "wave trough standard deviation Claus brightness temperature" ;
		stdctb:units = "K" ;
		stdctb:coordinates = "time lat lon" ;
		stdctb:cell_methods = "area: standard_deviation (over the wave trough)" ;
		stdctb:references = "Environmental Systems Science Centre (ESSC), [Robinson, G.J.] . Cloud Archive User Service (CLAUS), [Internet]. NCAS British Atmospheric Data Centre, 2002. Available from http://badc.nerc.ac.uk/view/badc.nerc.ac.uk__ATOM__dataent_claus." ;
	float ctb_area_fraction(sample) ;
		ctb_area_fraction:_FillValue = -999.f ;
		ctb_area_fraction:long_name = "wave trough Claus brightness temperature area fraction" ;
		ctb_area_fraction:units = "" ;
		ctb_area_fraction:coordinates = "time lat lon" ;
		ctb_area_fraction:references = "Environmental Systems Science Centre (ESSC), [Robinson, G.J.] . Cloud Archive User Service (CLAUS), [Internet]. NCAS British Atmospheric Data Centre, 2002. Available from http://badc.nerc.ac.uk/view/badc.nerc.ac.uk__ATOM__dataent_claus." ;
		ctb_area_fraction:comment = "Fractional area coverage of available Claus brightness temperature data for the wave trough." ;
	float meantpw(sample) ;
		meantpw:_FillValue = -999.f ;
		meantpw:long_name = "wave trough mean total precipitable water" ;
		meantpw:units = "mm" ;
		meantpw:coordinates = "time lat lon" ;
		meantpw:cell_methods = "area: mean (over the wave trough)" ;
		meantpw:platform = "DMSP SSM/I" ;
		meantpw:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		meantpw:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		meantpw:comment = "Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float stdtpw(sample) ;
		stdtpw:_FillValue = -999.f ;
		stdtpw:long_name = "wave trough standard deviation total precipitable water" ;
		stdtpw:units = "mm" ;
		stdtpw:coordinates = "time lat lon" ;
		stdtpw:cell_methods = "area: standard_deviation (over the wave trough)" ;
		stdtpw:platform = "DMSP SSM/I" ;
		stdtpw:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		stdtpw:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		stdtpw:comment = "Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float tpw_area_fraction(sample) ;
		tpw_area_fraction:_FillValue = -999.f ;
		tpw_area_fraction:long_name = "wave trough total precipitable water area fraction" ;
		tpw_area_fraction:coordinates = "time lat lon" ;
		tpw_area_fraction:platform = "DMSP SSM/I" ;
		tpw_area_fraction:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		tpw_area_fraction:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		tpw_area_fraction:comment = "Fractional area coverage of available SSM/I total precipitable water data for the wave trough. Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float meanrain(sample) ;
		meanrain:_FillValue = -999.f ;
		meanrain:long_name = "wave trough mean rain rate" ;
		meanrain:units = "mm hr-1" ;
		meanrain:coordinates = "time lat lon" ;
		meanrain:cell_methods = "area: mean (over the wave trough)" ;
		meanrain:platform = "DMSP SSM/I" ;
		meanrain:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		meanrain:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		meanrain:comment = "Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float stdrain(sample) ;
		stdrain:_FillValue = -999.f ;
		stdrain:long_name = "wave trough standard deviation rain rate" ;
		stdrain:units = "mm hr-1" ;
		stdrain:coordinates = "time lat lon" ;
		stdrain:cell_methods = "area: standard_deviation (over the wave trough)" ;
		stdrain:platform = "DMSP SSM/I" ;
		stdrain:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		stdrain:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		stdrain:comment = "Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float rain_area_fraction(sample) ;
		rain_area_fraction:_FillValue = -999.f ;
		rain_area_fraction:long_name = "wave trough total rain rate area fraction" ;
		rain_area_fraction:coordinates = "time lat lon" ;
		rain_area_fraction:platform = "DMSP SSM/I" ;
		rain_area_fraction:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		rain_area_fraction:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		rain_area_fraction:comment = "Fractional area coverage of available SSM/I rain rate data for the wave trough. Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float meancloud(sample) ;
		meancloud:_FillValue = -999.f ;
		meancloud:long_name = "wave trough mean total cloud liquid water" ;
		meancloud:units = "mm" ;
		meancloud:coordinates = "time lat lon" ;
		meancloud:cell_methods = "area: mean (over the wave trough)" ;
		meancloud:platform = "DMSP SSM/I" ;
		meancloud:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		meancloud:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		meancloud:comment = "Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float stdcloud(sample) ;
		stdcloud:_FillValue = -999.f ;
		stdcloud:long_name = "wave trough standard deviation cloud liquid water" ;
		stdcloud:units = "mm" ;
		stdcloud:coordinates = "time lat lon" ;
		stdcloud:cell_methods = "area: standard_deviation (over the wave trough)" ;
		stdcloud:platform = "DMSP SSM/I" ;
		stdcloud:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		stdcloud:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		stdcloud:comment = "Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;
	float cloud_area_fraction(sample) ;
		cloud_area_fraction:_FillValue = -999.f ;
		cloud_area_fraction:long_name = "wave trough total cloud liquid water area fraction" ;
		cloud_area_fraction:coordinates = "time lat lon" ;
		cloud_area_fraction:platform = "DMSP SSM/I" ;
		cloud_area_fraction:instrument = "F08:1987-1991, F10:1990-1997, F11:1991-2000, F13:1995-2009, F14:1997-2008, F15:1999-2006, F16:2003-2010, F17:2006-2010" ;
		cloud_area_fraction:references = "SSM/I and SSMIS data are produced by Remote Sensing Systems and sponsored by the NASA Earth Science MEaSUREs Program and are available at www.remss.com." ;
		cloud_area_fraction:comment = "Fractional area coverage of available SSM/I rain rate data for the wave trough. Satellite overpass data rounded to nearest 6-hr and averaged for all overlapping times and locations." ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:standard_name_vocabulary = "CF Standard Name Table (v26, 08 November 2013)" ;
		:title = "African Easterly Wave Climatology" ;
		:summary = "easterly wave trajectories for 700 hPa originating from Africa for 1987" ;
		:source = "NCEP Climate Forecast System Reanalysis" ;
		:id = "CFS_ew_700hPa_1987_AFR.nc" ;
		:naming_authority = "gov.noaa.ncdc" ;
		:time_coverage_start = "1987-01-01T00:00:00Z" ;
		:time_coverage_end = "1987-12-31T18:00:00Z" ;
		:time_coverage_resolution = "P6H" ;
		:time_coverage_duration = "P1Y" ;
		:geospatial_lat_min = -35.f ;
		:geospatial_lat_max = 35.f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = -140.f ;
		:geospatial_lon_max = 40.f ;
		:geospatial_lon_units = "degrees_north" ;
		:institution = "GATECH/GTRI > Georgia Institute of Technology, Georgia Tech Research Institute, School of Earth & Atmospheric Sciences" ;
		:creator_name = "James Belanger, Mark Jelinek, Judith Curry" ;
		:creator_email = "james.belanger@gatech.edu" ;
		:project = "U.S. Department of Commerce NOAA Grant 3506G58; National Science Foundation Grant 3506G42" ;
		:processing_level = "Level 4" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Earth Science Keywords, Version 8.0" ;
		:keywords = "EARTH SCIENCE, ATMOSPHERE, ATMOSPHERIC PHENOMENA, HURRICANES" ;
		:references = "Belanger, J.I, M. T. Jelinek, and  J. A. Curry, 2014: Revisiting the tropical cyclone-easterly wave relationship on interannual time scales, J. Climate." ;
		:date_created = "2014-07-25" ;
		:license = "No constraints on data access or use" ;
		:metadata_link = "gov.noaa.ncdc:C00784" ;
}
