netcdf tmpcdltest {
variables:
        int gfsmos_process_chain;
        gfsmos_process_chain:OM_Process = "(step1 step2)";

int step1;
        step1:LE_ProcessStep = "https://codes.nws.noaa.gov/NumericalWeatherPrediction/Models/GFS13" ;
        step1:LE_Source = "https://codes.nws.noaa.gov/DataAssimilation/Methods/GDAS13" ;

int step2;
        step2:LE_ProcessStep = "https://codes.nws.noaa.gov/StatisticalPostProcessing/Methods/GFSMOS05" ;
        step2:LE_Source = "https://codes.nws.noaa.gov/NumericalWeatherPrediction/Models/GFS13" ;

//global attribute
        :process_chain = "gfsmos_process_chain";
}
